This is an RTL file
this is a new line added from ws1
