This is a Testbench file in systemverilog
