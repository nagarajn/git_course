This is an RTL file
This can be another line in the rtl
this is a new line added from ws1
