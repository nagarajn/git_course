This is an RTL file
This can be another line in the rtl
