This is an RTL file
